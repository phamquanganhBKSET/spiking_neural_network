`define DATA_WIDTH   32                    // Buffer data width
`define BUFFER_DEPTH 4                     // Buffer depth
`define BUFFER_WIDTH $clog2(`BUFFER_DEPTH) // Buffer width
`define NUM_AXON     256                   // Number of axons
`define NUM_NEURON   256                   // Number of neurons
`define PACKET_WIDTH 30                    // Packet width
`define DX_MSB       29
`define DX_LSB       21
`define DY_MSB       20
`define DY_LSB       12
`define EAST         1
